module main

import list_utils

fn main() {
	println('Hello World!')
}
